library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity OSDBoot_832_ROM is
generic
	(
		maxAddrBitBRAM : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(maxAddrBitBRAM-2 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111";
	-- Second port
	addr2 : in std_logic_vector(maxAddrBitBRAM-2 downto 0) := (others=>'0');
	q2 : out std_logic_vector(31 downto 0);
	d2 : in std_logic_vector(31 downto 0) := X"00000000";
	we2 : in std_logic := '0';
	bytesel2 : in std_logic_vector(3 downto 0) := "1111"	
);
end OSDBoot_832_ROM;

architecture arch of OSDBoot_832_ROM is

type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
type ram_type is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

signal ram : ram_type :=
(
     0 => (x"01",x"da",x"87",x"04"),
     1 => (x"dd",x"87",x"0e",x"58"),
     2 => (x"5e",x"59",x"5a",x"0e"),
     3 => (x"27",x"00",x"00",x"00"),
     4 => (x"29",x"0f",x"26",x"4a"),
     5 => (x"26",x"49",x"26",x"48"),
     6 => (x"ff",x"80",x"26",x"08"),
     7 => (x"4f",x"27",x"00",x"00"),
     8 => (x"00",x"2d",x"4f",x"27"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"4f",x"4f",x"00",x"fd"),
    11 => (x"87",x"c1",x"ca",x"e0"),
    12 => (x"4e",x"c9",x"c0",x"48"),
    13 => (x"c2",x"28",x"c1",x"d5"),
    14 => (x"ea",x"e5",x"d6",x"ea"),
    15 => (x"49",x"71",x"46",x"c1"),
    16 => (x"88",x"01",x"f9",x"87"),
    17 => (x"c1",x"ca",x"e0",x"49"),
    18 => (x"c1",x"c1",x"cc",x"48"),
    19 => (x"89",x"d0",x"89",x"03"),
    20 => (x"c0",x"40",x"40",x"40"),
    21 => (x"40",x"f6",x"87",x"d0"),
    22 => (x"81",x"05",x"c0",x"50"),
    23 => (x"c1",x"89",x"05",x"f9"),
    24 => (x"87",x"c1",x"c1",x"ca"),
    25 => (x"4d",x"c1",x"c1",x"ca"),
    26 => (x"4c",x"74",x"ad",x"02"),
    27 => (x"c4",x"87",x"24",x"0f"),
    28 => (x"f7",x"87",x"c2",x"dc"),
    29 => (x"87",x"c1",x"c1",x"ca"),
    30 => (x"4d",x"c1",x"c1",x"ca"),
    31 => (x"4c",x"74",x"ad",x"02"),
    32 => (x"c6",x"87",x"c4",x"8c"),
    33 => (x"6c",x"0f",x"f5",x"87"),
    34 => (x"00",x"98",x"fc",x"87"),
    35 => (x"0e",x"5e",x"5b",x"5c"),
    36 => (x"0e",x"c4",x"c0",x"c0"),
    37 => (x"c0",x"4b",x"c9",x"d0"),
    38 => (x"4c",x"c9",x"e2",x"bf"),
    39 => (x"4a",x"49",x"c1",x"8a"),
    40 => (x"71",x"99",x"02",x"cf"),
    41 => (x"87",x"74",x"49",x"c1"),
    42 => (x"84",x"11",x"53",x"72"),
    43 => (x"49",x"c1",x"8a",x"71"),
    44 => (x"99",x"05",x"f1",x"87"),
    45 => (x"c2",x"87",x"26",x"4d"),
    46 => (x"26",x"4c",x"26",x"4b"),
    47 => (x"26",x"4f",x"1e",x"73"),
    48 => (x"1e",x"71",x"4b",x"e7"),
    49 => (x"48",x"c0",x"e0",x"50"),
    50 => (x"e3",x"48",x"c8",x"50"),
    51 => (x"e3",x"48",x"c6",x"50"),
    52 => (x"e7",x"48",x"c0",x"e1"),
    53 => (x"50",x"73",x"4a",x"c8"),
    54 => (x"b7",x"2a",x"c4",x"c0"),
    55 => (x"c0",x"c0",x"49",x"ca"),
    56 => (x"81",x"72",x"51",x"73"),
    57 => (x"4a",x"c3",x"ff",x"9a"),
    58 => (x"c4",x"c0",x"c0",x"c0"),
    59 => (x"49",x"cb",x"81",x"72"),
    60 => (x"51",x"e7",x"48",x"c0"),
    61 => (x"e0",x"50",x"e3",x"48"),
    62 => (x"c8",x"50",x"e3",x"48"),
    63 => (x"c0",x"50",x"e7",x"48"),
    64 => (x"c0",x"e1",x"50",x"fe"),
    65 => (x"f4",x"87",x"1e",x"73"),
    66 => (x"1e",x"c2",x"c0",x"c0"),
    67 => (x"4b",x"0f",x"fe",x"e9"),
    68 => (x"87",x"1e",x"73",x"1e"),
    69 => (x"eb",x"48",x"c3",x"ef"),
    70 => (x"50",x"e7",x"48",x"c0"),
    71 => (x"e0",x"50",x"e3",x"48"),
    72 => (x"c8",x"50",x"e3",x"48"),
    73 => (x"c6",x"50",x"e7",x"48"),
    74 => (x"c0",x"e1",x"50",x"ff"),
    75 => (x"c2",x"48",x"c1",x"9f"),
    76 => (x"78",x"e7",x"48",x"c0"),
    77 => (x"e0",x"50",x"e3",x"48"),
    78 => (x"c4",x"50",x"e3",x"48"),
    79 => (x"c2",x"50",x"e7",x"48"),
    80 => (x"c0",x"e1",x"50",x"e7"),
    81 => (x"48",x"c0",x"e0",x"50"),
    82 => (x"e3",x"48",x"c8",x"50"),
    83 => (x"e3",x"48",x"c7",x"50"),
    84 => (x"e7",x"48",x"c0",x"e1"),
    85 => (x"50",x"fc",x"f4",x"87"),
    86 => (x"c0",x"ff",x"ff",x"49"),
    87 => (x"fd",x"df",x"87",x"c0"),
    88 => (x"fc",x"c0",x"4b",x"c8"),
    89 => (x"dc",x"49",x"c0",x"f9"),
    90 => (x"d7",x"87",x"cd",x"e5"),
    91 => (x"87",x"70",x"98",x"02"),
    92 => (x"c1",x"c3",x"87",x"c0"),
    93 => (x"ff",x"f0",x"4b",x"c8"),
    94 => (x"c5",x"49",x"c0",x"f9"),
    95 => (x"c3",x"87",x"d3",x"cf"),
    96 => (x"87",x"70",x"98",x"02"),
    97 => (x"c0",x"e6",x"87",x"c3"),
    98 => (x"f0",x"4b",x"c2",x"c0"),
    99 => (x"c0",x"1e",x"c7",x"c8"),
   100 => (x"49",x"c0",x"ea",x"ef"),
   101 => (x"87",x"c4",x"86",x"70"),
   102 => (x"98",x"02",x"c8",x"87"),
   103 => (x"c3",x"ff",x"4b",x"fd"),
   104 => (x"e4",x"87",x"d9",x"87"),
   105 => (x"c7",x"d4",x"49",x"c0"),
   106 => (x"f8",x"d6",x"87",x"d0"),
   107 => (x"87",x"c7",x"e9",x"49"),
   108 => (x"c0",x"f8",x"cd",x"87"),
   109 => (x"c7",x"87",x"c8",x"f2"),
   110 => (x"49",x"c0",x"f8",x"c4"),
   111 => (x"87",x"73",x"49",x"fb"),
   112 => (x"fc",x"87",x"fe",x"da"),
   113 => (x"87",x"fb",x"f2",x"87"),
   114 => (x"38",x"33",x"32",x"4f"),
   115 => (x"53",x"44",x"41",x"44"),
   116 => (x"42",x"49",x"4e",x"00"),
   117 => (x"43",x"61",x"6e",x"27"),
   118 => (x"74",x"20",x"6c",x"6f"),
   119 => (x"61",x"64",x"20",x"66"),
   120 => (x"69",x"72",x"6d",x"77"),
   121 => (x"61",x"72",x"65",x"0a"),
   122 => (x"00",x"55",x"6e",x"61"),
   123 => (x"62",x"6c",x"65",x"20"),
   124 => (x"74",x"6f",x"20",x"6c"),
   125 => (x"6f",x"63",x"61",x"74"),
   126 => (x"65",x"20",x"70",x"61"),
   127 => (x"72",x"74",x"69",x"74"),
   128 => (x"69",x"6f",x"6e",x"0a"),
   129 => (x"00",x"48",x"75",x"6e"),
   130 => (x"74",x"69",x"6e",x"67"),
   131 => (x"20",x"66",x"6f",x"72"),
   132 => (x"20",x"70",x"61",x"72"),
   133 => (x"74",x"69",x"74",x"69"),
   134 => (x"6f",x"6e",x"0a",x"00"),
   135 => (x"49",x"6e",x"69",x"74"),
   136 => (x"69",x"61",x"6c",x"69"),
   137 => (x"7a",x"69",x"6e",x"67"),
   138 => (x"20",x"53",x"44",x"20"),
   139 => (x"63",x"61",x"72",x"64"),
   140 => (x"0a",x"00",x"46",x"61"),
   141 => (x"69",x"6c",x"65",x"64"),
   142 => (x"20",x"74",x"6f",x"20"),
   143 => (x"69",x"6e",x"69",x"74"),
   144 => (x"69",x"61",x"6c",x"69"),
   145 => (x"7a",x"65",x"20",x"53"),
   146 => (x"44",x"20",x"63",x"61"),
   147 => (x"72",x"64",x"0a",x"00"),
   148 => (x"00",x"00",x"00",x"00"),
   149 => (x"00",x"00",x"00",x"08"),
   150 => (x"33",x"fc",x"0f",x"ff"),
   151 => (x"00",x"df",x"f1",x"80"),
   152 => (x"60",x"f6",x"00",x"00"),
   153 => (x"00",x"12",x"1e",x"e4"),
   154 => (x"86",x"e3",x"48",x"c3"),
   155 => (x"ff",x"50",x"e3",x"97"),
   156 => (x"bf",x"7e",x"6e",x"49"),
   157 => (x"c3",x"ff",x"99",x"e3"),
   158 => (x"48",x"c3",x"ff",x"50"),
   159 => (x"c8",x"31",x"e3",x"97"),
   160 => (x"bf",x"48",x"c8",x"a6"),
   161 => (x"58",x"c3",x"ff",x"98"),
   162 => (x"cc",x"a6",x"58",x"70"),
   163 => (x"b1",x"e3",x"48",x"c3"),
   164 => (x"ff",x"50",x"c8",x"31"),
   165 => (x"e3",x"97",x"bf",x"48"),
   166 => (x"d0",x"a6",x"58",x"c3"),
   167 => (x"ff",x"98",x"d4",x"a6"),
   168 => (x"58",x"70",x"b1",x"e3"),
   169 => (x"48",x"c3",x"ff",x"50"),
   170 => (x"c8",x"31",x"e3",x"97"),
   171 => (x"bf",x"48",x"d8",x"a6"),
   172 => (x"58",x"c3",x"ff",x"98"),
   173 => (x"dc",x"a6",x"58",x"70"),
   174 => (x"b1",x"71",x"48",x"e4"),
   175 => (x"8e",x"26",x"4f",x"0e"),
   176 => (x"5e",x"5b",x"5c",x"0e"),
   177 => (x"1e",x"71",x"4a",x"49"),
   178 => (x"c3",x"ff",x"99",x"e3"),
   179 => (x"48",x"71",x"50",x"c1"),
   180 => (x"c1",x"cc",x"bf",x"05"),
   181 => (x"c8",x"87",x"d0",x"66"),
   182 => (x"48",x"c9",x"30",x"d4"),
   183 => (x"a6",x"58",x"d0",x"66"),
   184 => (x"49",x"d8",x"29",x"c3"),
   185 => (x"ff",x"99",x"e3",x"48"),
   186 => (x"71",x"50",x"d0",x"66"),
   187 => (x"49",x"d0",x"29",x"c3"),
   188 => (x"ff",x"99",x"e3",x"48"),
   189 => (x"71",x"50",x"d0",x"66"),
   190 => (x"49",x"c8",x"29",x"c3"),
   191 => (x"ff",x"99",x"e3",x"48"),
   192 => (x"71",x"50",x"d0",x"66"),
   193 => (x"49",x"c3",x"ff",x"99"),
   194 => (x"e3",x"48",x"71",x"50"),
   195 => (x"72",x"49",x"d0",x"29"),
   196 => (x"c3",x"ff",x"99",x"e3"),
   197 => (x"48",x"71",x"50",x"e3"),
   198 => (x"97",x"bf",x"7e",x"6e"),
   199 => (x"4b",x"c3",x"ff",x"9b"),
   200 => (x"c9",x"f0",x"ff",x"4c"),
   201 => (x"c3",x"ff",x"ab",x"05"),
   202 => (x"d9",x"87",x"e3",x"48"),
   203 => (x"c3",x"ff",x"50",x"e3"),
   204 => (x"97",x"bf",x"7e",x"6e"),
   205 => (x"4b",x"c3",x"ff",x"9b"),
   206 => (x"c1",x"8c",x"02",x"c6"),
   207 => (x"87",x"c3",x"ff",x"ab"),
   208 => (x"02",x"e7",x"87",x"73"),
   209 => (x"4a",x"c4",x"b7",x"2a"),
   210 => (x"c0",x"f0",x"a2",x"49"),
   211 => (x"c0",x"e6",x"ec",x"87"),
   212 => (x"73",x"4a",x"cf",x"9a"),
   213 => (x"c0",x"f0",x"a2",x"49"),
   214 => (x"c0",x"e6",x"e0",x"87"),
   215 => (x"73",x"48",x"26",x"c2"),
   216 => (x"87",x"26",x"4d",x"26"),
   217 => (x"4c",x"26",x"4b",x"26"),
   218 => (x"4f",x"1e",x"c0",x"49"),
   219 => (x"e3",x"48",x"c3",x"ff"),
   220 => (x"50",x"c1",x"81",x"c3"),
   221 => (x"c8",x"b7",x"a9",x"04"),
   222 => (x"f2",x"87",x"26",x"4f"),
   223 => (x"1e",x"73",x"1e",x"e8"),
   224 => (x"87",x"c4",x"f8",x"df"),
   225 => (x"4b",x"c0",x"1e",x"c0"),
   226 => (x"ff",x"f0",x"c1",x"f7"),
   227 => (x"49",x"fc",x"ef",x"87"),
   228 => (x"c4",x"86",x"c1",x"a8"),
   229 => (x"05",x"c0",x"e8",x"87"),
   230 => (x"e3",x"48",x"c3",x"ff"),
   231 => (x"50",x"c1",x"c0",x"c0"),
   232 => (x"c0",x"c0",x"c0",x"1e"),
   233 => (x"c0",x"e1",x"f0",x"c1"),
   234 => (x"e9",x"49",x"fc",x"d2"),
   235 => (x"87",x"c4",x"86",x"70"),
   236 => (x"98",x"05",x"c9",x"87"),
   237 => (x"e3",x"48",x"c3",x"ff"),
   238 => (x"50",x"c1",x"48",x"cb"),
   239 => (x"87",x"fe",x"e9",x"87"),
   240 => (x"c1",x"8b",x"05",x"fe"),
   241 => (x"ff",x"87",x"c0",x"48"),
   242 => (x"fe",x"da",x"87",x"1e"),
   243 => (x"73",x"1e",x"e3",x"48"),
   244 => (x"c3",x"ff",x"50",x"d0"),
   245 => (x"c5",x"49",x"c0",x"ef"),
   246 => (x"e7",x"87",x"d3",x"4b"),
   247 => (x"c0",x"1e",x"c0",x"ff"),
   248 => (x"f0",x"c1",x"c1",x"49"),
   249 => (x"fb",x"d8",x"87",x"c4"),
   250 => (x"86",x"70",x"98",x"05"),
   251 => (x"c9",x"87",x"e3",x"48"),
   252 => (x"c3",x"ff",x"50",x"c1"),
   253 => (x"48",x"cb",x"87",x"fd"),
   254 => (x"ef",x"87",x"c1",x"8b"),
   255 => (x"05",x"ff",x"dc",x"87"),
   256 => (x"c0",x"48",x"fd",x"e0"),
   257 => (x"87",x"43",x"6d",x"64"),
   258 => (x"5f",x"69",x"6e",x"69"),
   259 => (x"74",x"0a",x"00",x"1e"),
   260 => (x"73",x"1e",x"1e",x"fd"),
   261 => (x"d3",x"87",x"c6",x"ea"),
   262 => (x"1e",x"c0",x"e1",x"f0"),
   263 => (x"c1",x"c8",x"49",x"fa"),
   264 => (x"dd",x"87",x"70",x"4b"),
   265 => (x"1e",x"d2",x"fb",x"1e"),
   266 => (x"c0",x"ee",x"c1",x"87"),
   267 => (x"cc",x"86",x"c1",x"ab"),
   268 => (x"02",x"c8",x"87",x"fe"),
   269 => (x"d5",x"87",x"c0",x"48"),
   270 => (x"c1",x"fc",x"87",x"f8"),
   271 => (x"e8",x"87",x"70",x"49"),
   272 => (x"cf",x"ff",x"ff",x"99"),
   273 => (x"c6",x"ea",x"a9",x"02"),
   274 => (x"c8",x"87",x"fd",x"fe"),
   275 => (x"87",x"c0",x"48",x"c1"),
   276 => (x"e5",x"87",x"e3",x"48"),
   277 => (x"c3",x"ff",x"50",x"c0"),
   278 => (x"f1",x"4b",x"fc",x"df"),
   279 => (x"87",x"70",x"98",x"02"),
   280 => (x"c1",x"c3",x"87",x"c0"),
   281 => (x"1e",x"c0",x"ff",x"f0"),
   282 => (x"c1",x"fa",x"49",x"f9"),
   283 => (x"d1",x"87",x"c4",x"86"),
   284 => (x"70",x"98",x"05",x"c0"),
   285 => (x"f0",x"87",x"e3",x"48"),
   286 => (x"c3",x"ff",x"50",x"e3"),
   287 => (x"97",x"bf",x"7e",x"6e"),
   288 => (x"49",x"c3",x"ff",x"99"),
   289 => (x"e3",x"48",x"c3",x"ff"),
   290 => (x"50",x"e3",x"48",x"c3"),
   291 => (x"ff",x"50",x"e3",x"48"),
   292 => (x"c3",x"ff",x"50",x"e3"),
   293 => (x"48",x"c3",x"ff",x"50"),
   294 => (x"c1",x"c0",x"99",x"02"),
   295 => (x"c4",x"87",x"c1",x"48"),
   296 => (x"d5",x"87",x"c0",x"48"),
   297 => (x"d1",x"87",x"c2",x"ab"),
   298 => (x"05",x"c4",x"87",x"c0"),
   299 => (x"48",x"c8",x"87",x"c1"),
   300 => (x"8b",x"05",x"fe",x"e5"),
   301 => (x"87",x"c0",x"48",x"26"),
   302 => (x"fa",x"ea",x"87",x"63"),
   303 => (x"6d",x"64",x"5f",x"43"),
   304 => (x"4d",x"44",x"38",x"20"),
   305 => (x"72",x"65",x"73",x"70"),
   306 => (x"6f",x"6e",x"73",x"65"),
   307 => (x"3a",x"20",x"25",x"64"),
   308 => (x"0a",x"00",x"1e",x"73"),
   309 => (x"1e",x"c1",x"c1",x"cc"),
   310 => (x"48",x"c1",x"78",x"eb"),
   311 => (x"48",x"c3",x"ef",x"50"),
   312 => (x"c7",x"4b",x"e7",x"48"),
   313 => (x"c3",x"50",x"fa",x"c0"),
   314 => (x"87",x"e7",x"48",x"c2"),
   315 => (x"50",x"e3",x"48",x"c3"),
   316 => (x"ff",x"50",x"c0",x"1e"),
   317 => (x"c0",x"e5",x"d0",x"c1"),
   318 => (x"c0",x"49",x"f7",x"c2"),
   319 => (x"87",x"c4",x"86",x"c1"),
   320 => (x"a8",x"05",x"c1",x"87"),
   321 => (x"4b",x"c2",x"ab",x"05"),
   322 => (x"c5",x"87",x"c0",x"48"),
   323 => (x"c0",x"ef",x"87",x"c1"),
   324 => (x"8b",x"05",x"ff",x"cd"),
   325 => (x"87",x"fb",x"f7",x"87"),
   326 => (x"c1",x"c1",x"d0",x"58"),
   327 => (x"70",x"98",x"05",x"cd"),
   328 => (x"87",x"c1",x"1e",x"c0"),
   329 => (x"ff",x"f0",x"c1",x"d0"),
   330 => (x"49",x"f6",x"d3",x"87"),
   331 => (x"c4",x"86",x"e3",x"48"),
   332 => (x"c3",x"ff",x"50",x"e7"),
   333 => (x"48",x"c3",x"50",x"e3"),
   334 => (x"48",x"c3",x"ff",x"50"),
   335 => (x"c1",x"48",x"f8",x"e4"),
   336 => (x"87",x"0e",x"5e",x"5b"),
   337 => (x"5c",x"5d",x"0e",x"1e"),
   338 => (x"71",x"4a",x"c0",x"4d"),
   339 => (x"e3",x"48",x"c3",x"ff"),
   340 => (x"50",x"e7",x"48",x"c2"),
   341 => (x"50",x"eb",x"48",x"c7"),
   342 => (x"50",x"e3",x"48",x"c3"),
   343 => (x"ff",x"50",x"72",x"1e"),
   344 => (x"c0",x"ff",x"f0",x"c1"),
   345 => (x"d1",x"49",x"f5",x"d6"),
   346 => (x"87",x"c4",x"86",x"70"),
   347 => (x"98",x"05",x"c1",x"c5"),
   348 => (x"87",x"c5",x"ee",x"cd"),
   349 => (x"df",x"4b",x"e3",x"48"),
   350 => (x"c3",x"ff",x"50",x"e3"),
   351 => (x"97",x"bf",x"7e",x"6e"),
   352 => (x"49",x"c3",x"ff",x"99"),
   353 => (x"c3",x"fe",x"a9",x"05"),
   354 => (x"dd",x"87",x"c0",x"4c"),
   355 => (x"f3",x"d7",x"87",x"d4"),
   356 => (x"66",x"08",x"78",x"d4"),
   357 => (x"66",x"48",x"c4",x"80"),
   358 => (x"d8",x"a6",x"58",x"c1"),
   359 => (x"84",x"c2",x"c0",x"b7"),
   360 => (x"ac",x"04",x"e8",x"87"),
   361 => (x"c1",x"4b",x"4d",x"c1"),
   362 => (x"8b",x"05",x"ff",x"c9"),
   363 => (x"87",x"e3",x"48",x"c3"),
   364 => (x"ff",x"50",x"e7",x"48"),
   365 => (x"c3",x"50",x"75",x"48"),
   366 => (x"26",x"f6",x"e5",x"87"),
   367 => (x"1e",x"73",x"1e",x"71"),
   368 => (x"4b",x"49",x"d8",x"29"),
   369 => (x"c3",x"ff",x"99",x"73"),
   370 => (x"4a",x"c8",x"2a",x"cf"),
   371 => (x"fc",x"c0",x"9a",x"72"),
   372 => (x"b1",x"73",x"4a",x"c8"),
   373 => (x"32",x"c0",x"ff",x"f0"),
   374 => (x"c0",x"c0",x"9a",x"72"),
   375 => (x"b1",x"73",x"4a",x"d8"),
   376 => (x"32",x"ff",x"c0",x"c0"),
   377 => (x"c0",x"c0",x"9a",x"72"),
   378 => (x"b1",x"71",x"48",x"c4"),
   379 => (x"87",x"26",x"4d",x"26"),
   380 => (x"4c",x"26",x"4b",x"26"),
   381 => (x"4f",x"1e",x"73",x"1e"),
   382 => (x"71",x"4b",x"49",x"c8"),
   383 => (x"29",x"c3",x"ff",x"99"),
   384 => (x"73",x"4a",x"c8",x"32"),
   385 => (x"cf",x"fc",x"c0",x"9a"),
   386 => (x"72",x"b1",x"71",x"48"),
   387 => (x"e3",x"87",x"0e",x"5e"),
   388 => (x"5b",x"5c",x"0e",x"71"),
   389 => (x"4b",x"c0",x"4c",x"d0"),
   390 => (x"66",x"48",x"c0",x"b7"),
   391 => (x"a8",x"06",x"c0",x"e3"),
   392 => (x"87",x"13",x"4a",x"cc"),
   393 => (x"66",x"97",x"bf",x"49"),
   394 => (x"cc",x"66",x"48",x"c1"),
   395 => (x"80",x"d0",x"a6",x"58"),
   396 => (x"71",x"b7",x"aa",x"02"),
   397 => (x"c4",x"87",x"c1",x"48"),
   398 => (x"cc",x"87",x"c1",x"84"),
   399 => (x"d0",x"66",x"b7",x"ac"),
   400 => (x"04",x"ff",x"dd",x"87"),
   401 => (x"c0",x"48",x"c2",x"87"),
   402 => (x"26",x"4d",x"26",x"4c"),
   403 => (x"26",x"4b",x"26",x"4f"),
   404 => (x"0e",x"5e",x"5b",x"5c"),
   405 => (x"0e",x"1e",x"c1",x"ca"),
   406 => (x"c0",x"48",x"ff",x"78"),
   407 => (x"c1",x"c9",x"d8",x"48"),
   408 => (x"c0",x"78",x"c0",x"e7"),
   409 => (x"c8",x"49",x"c0",x"e5"),
   410 => (x"d7",x"87",x"c1",x"c1"),
   411 => (x"d0",x"1e",x"c0",x"49"),
   412 => (x"fb",x"ce",x"87",x"c4"),
   413 => (x"86",x"70",x"98",x"05"),
   414 => (x"c5",x"87",x"c0",x"48"),
   415 => (x"cb",x"c2",x"87",x"c0"),
   416 => (x"4b",x"c1",x"c9",x"fc"),
   417 => (x"48",x"c1",x"78",x"c8"),
   418 => (x"1e",x"c0",x"e7",x"d5"),
   419 => (x"1e",x"c1",x"c2",x"c6"),
   420 => (x"49",x"fd",x"fa",x"87"),
   421 => (x"c8",x"86",x"70",x"98"),
   422 => (x"05",x"c6",x"87",x"c1"),
   423 => (x"c9",x"fc",x"48",x"c0"),
   424 => (x"78",x"c8",x"1e",x"c0"),
   425 => (x"e7",x"de",x"1e",x"c1"),
   426 => (x"c2",x"e2",x"49",x"fd"),
   427 => (x"e0",x"87",x"c8",x"86"),
   428 => (x"70",x"98",x"05",x"c6"),
   429 => (x"87",x"c1",x"c9",x"fc"),
   430 => (x"48",x"c0",x"78",x"c8"),
   431 => (x"1e",x"c0",x"e7",x"e7"),
   432 => (x"1e",x"c1",x"c2",x"e2"),
   433 => (x"49",x"fd",x"c6",x"87"),
   434 => (x"c8",x"86",x"70",x"98"),
   435 => (x"05",x"c5",x"87",x"c0"),
   436 => (x"48",x"c9",x"ed",x"87"),
   437 => (x"c1",x"c9",x"fc",x"bf"),
   438 => (x"1e",x"c0",x"e7",x"f0"),
   439 => (x"1e",x"c0",x"e3",x"cc"),
   440 => (x"87",x"c8",x"86",x"c1"),
   441 => (x"c9",x"fc",x"bf",x"02"),
   442 => (x"c1",x"ef",x"87",x"c1"),
   443 => (x"c1",x"d0",x"4a",x"48"),
   444 => (x"c6",x"fe",x"a0",x"4c"),
   445 => (x"c1",x"c8",x"d6",x"bf"),
   446 => (x"4b",x"c1",x"c9",x"ce"),
   447 => (x"9f",x"bf",x"49",x"72"),
   448 => (x"7e",x"c5",x"d6",x"ea"),
   449 => (x"a9",x"05",x"c0",x"cd"),
   450 => (x"87",x"c8",x"a4",x"4a"),
   451 => (x"6a",x"49",x"fa",x"eb"),
   452 => (x"87",x"70",x"49",x"4b"),
   453 => (x"dc",x"87",x"c7",x"fe"),
   454 => (x"a2",x"49",x"9f",x"69"),
   455 => (x"49",x"ca",x"e9",x"d5"),
   456 => (x"a9",x"02",x"c0",x"cd"),
   457 => (x"87",x"c0",x"e5",x"c5"),
   458 => (x"49",x"c0",x"e2",x"d4"),
   459 => (x"87",x"c0",x"48",x"c8"),
   460 => (x"cf",x"87",x"73",x"1e"),
   461 => (x"c0",x"e5",x"e3",x"1e"),
   462 => (x"c0",x"e1",x"f1",x"87"),
   463 => (x"c1",x"c1",x"d0",x"1e"),
   464 => (x"73",x"49",x"f7",x"fc"),
   465 => (x"87",x"cc",x"86",x"70"),
   466 => (x"98",x"05",x"c0",x"c5"),
   467 => (x"87",x"c0",x"48",x"c7"),
   468 => (x"ef",x"87",x"c0",x"e5"),
   469 => (x"fb",x"49",x"c0",x"e1"),
   470 => (x"e7",x"87",x"c0",x"e8"),
   471 => (x"c3",x"1e",x"c0",x"e1"),
   472 => (x"cb",x"87",x"c8",x"1e"),
   473 => (x"c0",x"e8",x"db",x"1e"),
   474 => (x"c1",x"c2",x"e2",x"49"),
   475 => (x"fa",x"df",x"87",x"cc"),
   476 => (x"86",x"70",x"98",x"05"),
   477 => (x"c0",x"c9",x"87",x"c1"),
   478 => (x"c9",x"d8",x"48",x"c1"),
   479 => (x"78",x"c0",x"e4",x"87"),
   480 => (x"c8",x"1e",x"c0",x"e8"),
   481 => (x"e4",x"1e",x"c1",x"c2"),
   482 => (x"c6",x"49",x"fa",x"c1"),
   483 => (x"87",x"c8",x"86",x"70"),
   484 => (x"98",x"02",x"c0",x"cf"),
   485 => (x"87",x"c0",x"e6",x"e2"),
   486 => (x"1e",x"c0",x"e0",x"d0"),
   487 => (x"87",x"c4",x"86",x"c0"),
   488 => (x"48",x"c6",x"dd",x"87"),
   489 => (x"c1",x"c9",x"ce",x"97"),
   490 => (x"bf",x"49",x"c1",x"d5"),
   491 => (x"a9",x"05",x"c0",x"cd"),
   492 => (x"87",x"c1",x"c9",x"cf"),
   493 => (x"97",x"bf",x"49",x"c2"),
   494 => (x"ea",x"a9",x"02",x"c0"),
   495 => (x"c5",x"87",x"c0",x"48"),
   496 => (x"c5",x"fe",x"87",x"c1"),
   497 => (x"c1",x"d0",x"97",x"bf"),
   498 => (x"49",x"c3",x"e9",x"a9"),
   499 => (x"02",x"c0",x"d2",x"87"),
   500 => (x"c1",x"c1",x"d0",x"97"),
   501 => (x"bf",x"49",x"c3",x"eb"),
   502 => (x"a9",x"02",x"c0",x"c5"),
   503 => (x"87",x"c0",x"48",x"c5"),
   504 => (x"df",x"87",x"c1",x"c1"),
   505 => (x"db",x"97",x"bf",x"49"),
   506 => (x"99",x"05",x"c0",x"cc"),
   507 => (x"87",x"c1",x"c1",x"dc"),
   508 => (x"97",x"bf",x"49",x"c2"),
   509 => (x"a9",x"02",x"c0",x"c5"),
   510 => (x"87",x"c0",x"48",x"c5"),
   511 => (x"c3",x"87",x"c1",x"c1"),
   512 => (x"dd",x"97",x"bf",x"48"),
   513 => (x"c1",x"c9",x"d4",x"58"),
   514 => (x"70",x"49",x"c1",x"89"),
   515 => (x"c1",x"c9",x"d8",x"59"),
   516 => (x"c1",x"c1",x"de",x"97"),
   517 => (x"bf",x"49",x"73",x"81"),
   518 => (x"c1",x"c1",x"df",x"97"),
   519 => (x"bf",x"4a",x"c8",x"32"),
   520 => (x"c1",x"c9",x"dc",x"48"),
   521 => (x"72",x"a1",x"78",x"c1"),
   522 => (x"c1",x"e0",x"97",x"bf"),
   523 => (x"48",x"c1",x"c9",x"f4"),
   524 => (x"58",x"c1",x"c9",x"d8"),
   525 => (x"bf",x"02",x"c2",x"ea"),
   526 => (x"87",x"c8",x"1e",x"c0"),
   527 => (x"e6",x"ff",x"1e",x"c1"),
   528 => (x"c2",x"e2",x"49",x"f7"),
   529 => (x"c8",x"87",x"c8",x"86"),
   530 => (x"70",x"98",x"02",x"c0"),
   531 => (x"c5",x"87",x"c0",x"48"),
   532 => (x"c3",x"ee",x"87",x"c1"),
   533 => (x"c9",x"d0",x"bf",x"48"),
   534 => (x"c4",x"30",x"c1",x"c9"),
   535 => (x"f8",x"58",x"c1",x"c9"),
   536 => (x"d0",x"bf",x"4a",x"c1"),
   537 => (x"c9",x"f0",x"5a",x"c1"),
   538 => (x"c1",x"f5",x"97",x"bf"),
   539 => (x"49",x"c8",x"31",x"c1"),
   540 => (x"c1",x"f4",x"97",x"bf"),
   541 => (x"4b",x"a1",x"49",x"c1"),
   542 => (x"c1",x"f6",x"97",x"bf"),
   543 => (x"4b",x"d0",x"33",x"73"),
   544 => (x"a1",x"49",x"c1",x"c1"),
   545 => (x"f7",x"97",x"bf",x"4b"),
   546 => (x"d8",x"33",x"73",x"a1"),
   547 => (x"49",x"c1",x"c9",x"fc"),
   548 => (x"59",x"c1",x"c9",x"f0"),
   549 => (x"bf",x"49",x"c1",x"c9"),
   550 => (x"f8",x"bf",x"91",x"c1"),
   551 => (x"c9",x"dc",x"bf",x"81"),
   552 => (x"c1",x"c9",x"e4",x"59"),
   553 => (x"c1",x"c1",x"fd",x"97"),
   554 => (x"bf",x"4b",x"c8",x"33"),
   555 => (x"c1",x"c1",x"fc",x"97"),
   556 => (x"bf",x"4c",x"a3",x"4b"),
   557 => (x"c1",x"c1",x"fe",x"97"),
   558 => (x"bf",x"4c",x"d0",x"34"),
   559 => (x"74",x"a3",x"4b",x"c1"),
   560 => (x"c1",x"ff",x"97",x"bf"),
   561 => (x"4c",x"cf",x"9c",x"d8"),
   562 => (x"34",x"74",x"a3",x"4b"),
   563 => (x"c1",x"c9",x"e8",x"5b"),
   564 => (x"c1",x"c9",x"e4",x"bf"),
   565 => (x"4b",x"c2",x"8b",x"73"),
   566 => (x"92",x"c1",x"c9",x"e8"),
   567 => (x"48",x"72",x"a1",x"78"),
   568 => (x"c1",x"dc",x"87",x"c1"),
   569 => (x"c1",x"e2",x"97",x"bf"),
   570 => (x"49",x"c8",x"31",x"c1"),
   571 => (x"c1",x"e1",x"97",x"bf"),
   572 => (x"4a",x"a1",x"49",x"c1"),
   573 => (x"c9",x"f8",x"59",x"c1"),
   574 => (x"c9",x"f4",x"bf",x"49"),
   575 => (x"c5",x"31",x"c7",x"ff"),
   576 => (x"81",x"c9",x"29",x"c1"),
   577 => (x"c9",x"f0",x"59",x"c1"),
   578 => (x"c1",x"e7",x"97",x"bf"),
   579 => (x"49",x"c8",x"31",x"c1"),
   580 => (x"c1",x"e6",x"97",x"bf"),
   581 => (x"4a",x"a1",x"49",x"c1"),
   582 => (x"c9",x"fc",x"59",x"c1"),
   583 => (x"c9",x"f0",x"bf",x"49"),
   584 => (x"c1",x"c9",x"f8",x"bf"),
   585 => (x"91",x"c1",x"c9",x"dc"),
   586 => (x"bf",x"81",x"c1",x"c9"),
   587 => (x"ec",x"59",x"c1",x"c9"),
   588 => (x"e4",x"48",x"c0",x"78"),
   589 => (x"c1",x"c9",x"ec",x"bf"),
   590 => (x"48",x"71",x"80",x"c1"),
   591 => (x"c9",x"e4",x"58",x"c1"),
   592 => (x"48",x"26",x"f4",x"c5"),
   593 => (x"87",x"4e",x"6f",x"20"),
   594 => (x"70",x"61",x"72",x"74"),
   595 => (x"69",x"74",x"69",x"6f"),
   596 => (x"6e",x"20",x"73",x"69"),
   597 => (x"67",x"6e",x"61",x"74"),
   598 => (x"75",x"72",x"65",x"20"),
   599 => (x"66",x"6f",x"75",x"6e"),
   600 => (x"64",x"0a",x"00",x"52"),
   601 => (x"65",x"61",x"64",x"69"),
   602 => (x"6e",x"67",x"20",x"62"),
   603 => (x"6f",x"6f",x"74",x"20"),
   604 => (x"73",x"65",x"63",x"74"),
   605 => (x"6f",x"72",x"20",x"25"),
   606 => (x"64",x"0a",x"00",x"52"),
   607 => (x"65",x"61",x"64",x"20"),
   608 => (x"62",x"6f",x"6f",x"74"),
   609 => (x"20",x"73",x"65",x"63"),
   610 => (x"74",x"6f",x"72",x"20"),
   611 => (x"66",x"72",x"6f",x"6d"),
   612 => (x"20",x"66",x"69",x"72"),
   613 => (x"73",x"74",x"20",x"70"),
   614 => (x"61",x"72",x"74",x"69"),
   615 => (x"74",x"69",x"6f",x"6e"),
   616 => (x"0a",x"00",x"55",x"6e"),
   617 => (x"73",x"75",x"70",x"70"),
   618 => (x"6f",x"72",x"74",x"65"),
   619 => (x"64",x"20",x"70",x"61"),
   620 => (x"72",x"74",x"69",x"74"),
   621 => (x"69",x"6f",x"6e",x"20"),
   622 => (x"74",x"79",x"70",x"65"),
   623 => (x"21",x"0d",x"00",x"46"),
   624 => (x"41",x"54",x"33",x"32"),
   625 => (x"20",x"20",x"20",x"00"),
   626 => (x"52",x"65",x"61",x"64"),
   627 => (x"69",x"6e",x"67",x"20"),
   628 => (x"4d",x"42",x"52",x"0a"),
   629 => (x"00",x"46",x"41",x"54"),
   630 => (x"31",x"36",x"20",x"20"),
   631 => (x"20",x"00",x"46",x"41"),
   632 => (x"54",x"33",x"32",x"20"),
   633 => (x"20",x"20",x"00",x"46"),
   634 => (x"41",x"54",x"31",x"32"),
   635 => (x"20",x"20",x"20",x"00"),
   636 => (x"50",x"61",x"72",x"74"),
   637 => (x"69",x"74",x"69",x"6f"),
   638 => (x"6e",x"63",x"6f",x"75"),
   639 => (x"6e",x"74",x"20",x"25"),
   640 => (x"64",x"0a",x"00",x"48"),
   641 => (x"75",x"6e",x"74",x"69"),
   642 => (x"6e",x"67",x"20",x"66"),
   643 => (x"6f",x"72",x"20",x"66"),
   644 => (x"69",x"6c",x"65",x"73"),
   645 => (x"79",x"73",x"74",x"65"),
   646 => (x"6d",x"0a",x"00",x"46"),
   647 => (x"41",x"54",x"33",x"32"),
   648 => (x"20",x"20",x"20",x"00"),
   649 => (x"46",x"41",x"54",x"31"),
   650 => (x"36",x"20",x"20",x"20"),
   651 => (x"00",x"0e",x"5e",x"5b"),
   652 => (x"5c",x"5d",x"0e",x"71"),
   653 => (x"4a",x"c1",x"c9",x"d8"),
   654 => (x"bf",x"02",x"cc",x"87"),
   655 => (x"72",x"4b",x"c7",x"b7"),
   656 => (x"2b",x"72",x"4c",x"c1"),
   657 => (x"ff",x"9c",x"ca",x"87"),
   658 => (x"72",x"4b",x"c8",x"b7"),
   659 => (x"2b",x"72",x"4c",x"c3"),
   660 => (x"ff",x"9c",x"73",x"49"),
   661 => (x"c1",x"ca",x"c0",x"bf"),
   662 => (x"a9",x"02",x"c0",x"e0"),
   663 => (x"87",x"c1",x"c1",x"d0"),
   664 => (x"1e",x"73",x"4a",x"c1"),
   665 => (x"c9",x"dc",x"bf",x"49"),
   666 => (x"72",x"81",x"eb",x"d4"),
   667 => (x"87",x"c4",x"86",x"70"),
   668 => (x"98",x"05",x"c5",x"87"),
   669 => (x"c0",x"48",x"c0",x"f5"),
   670 => (x"87",x"c1",x"ca",x"c4"),
   671 => (x"5b",x"c1",x"c9",x"d8"),
   672 => (x"bf",x"02",x"d8",x"87"),
   673 => (x"74",x"4a",x"c4",x"92"),
   674 => (x"c1",x"c1",x"d0",x"82"),
   675 => (x"6a",x"49",x"ec",x"eb"),
   676 => (x"87",x"70",x"49",x"4d"),
   677 => (x"cf",x"ff",x"ff",x"ff"),
   678 => (x"ff",x"9d",x"d0",x"87"),
   679 => (x"74",x"4a",x"c2",x"92"),
   680 => (x"c1",x"c1",x"d0",x"82"),
   681 => (x"9f",x"6a",x"49",x"ed"),
   682 => (x"cb",x"87",x"70",x"4d"),
   683 => (x"75",x"48",x"ee",x"d7"),
   684 => (x"87",x"0e",x"5e",x"5b"),
   685 => (x"5c",x"5d",x"0e",x"f4"),
   686 => (x"86",x"71",x"4c",x"c0"),
   687 => (x"4b",x"c1",x"ca",x"c0"),
   688 => (x"48",x"ff",x"78",x"c1"),
   689 => (x"c9",x"e4",x"bf",x"7e"),
   690 => (x"c1",x"c9",x"e8",x"bf"),
   691 => (x"4d",x"c1",x"c9",x"d8"),
   692 => (x"bf",x"02",x"cb",x"87"),
   693 => (x"c1",x"c9",x"d0",x"bf"),
   694 => (x"49",x"c4",x"31",x"71"),
   695 => (x"4a",x"c7",x"87",x"c1"),
   696 => (x"c9",x"ec",x"bf",x"4a"),
   697 => (x"c4",x"32",x"c8",x"a6"),
   698 => (x"5a",x"c8",x"a6",x"48"),
   699 => (x"c0",x"78",x"c4",x"66"),
   700 => (x"48",x"c0",x"a8",x"06"),
   701 => (x"c3",x"c6",x"87",x"c8"),
   702 => (x"66",x"49",x"cf",x"99"),
   703 => (x"05",x"dd",x"87",x"75"),
   704 => (x"1e",x"c0",x"ef",x"fe"),
   705 => (x"1e",x"d2",x"e5",x"87"),
   706 => (x"c1",x"c1",x"d0",x"1e"),
   707 => (x"75",x"49",x"c1",x"85"),
   708 => (x"71",x"e8",x"ed",x"87"),
   709 => (x"cc",x"86",x"c1",x"c1"),
   710 => (x"d0",x"4b",x"c3",x"87"),
   711 => (x"c0",x"e0",x"83",x"97"),
   712 => (x"6b",x"49",x"99",x"02"),
   713 => (x"c2",x"c4",x"87",x"97"),
   714 => (x"6b",x"49",x"c3",x"e5"),
   715 => (x"a9",x"02",x"c1",x"fa"),
   716 => (x"87",x"cb",x"a3",x"49"),
   717 => (x"97",x"69",x"49",x"d8"),
   718 => (x"99",x"05",x"c1",x"ee"),
   719 => (x"87",x"cb",x"1e",x"c0"),
   720 => (x"e0",x"66",x"1e",x"73"),
   721 => (x"49",x"eb",x"c6",x"87"),
   722 => (x"c8",x"86",x"70",x"98"),
   723 => (x"05",x"c1",x"db",x"87"),
   724 => (x"dc",x"a3",x"4a",x"6a"),
   725 => (x"49",x"e9",x"e4",x"87"),
   726 => (x"70",x"4a",x"c4",x"a4"),
   727 => (x"49",x"72",x"79",x"da"),
   728 => (x"a3",x"4a",x"9f",x"6a"),
   729 => (x"49",x"ea",x"cd",x"87"),
   730 => (x"70",x"7e",x"c1",x"c9"),
   731 => (x"d8",x"bf",x"02",x"d8"),
   732 => (x"87",x"d4",x"a3",x"4a"),
   733 => (x"9f",x"6a",x"49",x"e9"),
   734 => (x"fb",x"87",x"70",x"49"),
   735 => (x"c0",x"ff",x"ff",x"99"),
   736 => (x"71",x"48",x"d0",x"30"),
   737 => (x"c8",x"a6",x"58",x"c5"),
   738 => (x"87",x"c4",x"a6",x"48"),
   739 => (x"c0",x"78",x"c4",x"66"),
   740 => (x"4a",x"6e",x"82",x"c8"),
   741 => (x"a4",x"49",x"72",x"79"),
   742 => (x"c0",x"7c",x"dc",x"66"),
   743 => (x"1e",x"c0",x"f0",x"db"),
   744 => (x"1e",x"d0",x"c9",x"87"),
   745 => (x"c8",x"86",x"c1",x"48"),
   746 => (x"c1",x"ce",x"87",x"c8"),
   747 => (x"66",x"48",x"c1",x"80"),
   748 => (x"cc",x"a6",x"58",x"c8"),
   749 => (x"66",x"48",x"c4",x"66"),
   750 => (x"a8",x"04",x"fc",x"fa"),
   751 => (x"87",x"c1",x"c9",x"d8"),
   752 => (x"bf",x"02",x"c0",x"f2"),
   753 => (x"87",x"6e",x"49",x"f9"),
   754 => (x"e3",x"87",x"70",x"49"),
   755 => (x"7e",x"1e",x"c0",x"f0"),
   756 => (x"ec",x"1e",x"cf",x"d8"),
   757 => (x"87",x"c8",x"86",x"6e"),
   758 => (x"49",x"cf",x"ff",x"ff"),
   759 => (x"ff",x"f8",x"99",x"a9"),
   760 => (x"02",x"d4",x"87",x"6e"),
   761 => (x"49",x"c2",x"89",x"c1"),
   762 => (x"c9",x"d0",x"bf",x"4a"),
   763 => (x"91",x"c1",x"c9",x"e0"),
   764 => (x"bf",x"4d",x"71",x"85"),
   765 => (x"fb",x"f2",x"87",x"c0"),
   766 => (x"48",x"f4",x"8e",x"e9"),
   767 => (x"ca",x"87",x"52",x"65"),
   768 => (x"61",x"64",x"69",x"6e"),
   769 => (x"67",x"20",x"64",x"69"),
   770 => (x"72",x"65",x"63",x"74"),
   771 => (x"6f",x"72",x"79",x"20"),
   772 => (x"73",x"65",x"63",x"74"),
   773 => (x"6f",x"72",x"20",x"25"),
   774 => (x"64",x"0a",x"00",x"66"),
   775 => (x"69",x"6c",x"65",x"20"),
   776 => (x"22",x"25",x"73",x"22"),
   777 => (x"20",x"66",x"6f",x"75"),
   778 => (x"6e",x"64",x"0d",x"00"),
   779 => (x"47",x"65",x"74",x"46"),
   780 => (x"41",x"54",x"4c",x"69"),
   781 => (x"6e",x"6b",x"20",x"72"),
   782 => (x"65",x"74",x"75",x"72"),
   783 => (x"6e",x"65",x"64",x"20"),
   784 => (x"25",x"64",x"0a",x"00"),
   785 => (x"0e",x"5e",x"5b",x"5c"),
   786 => (x"5d",x"0e",x"1e",x"71"),
   787 => (x"4b",x"1e",x"c1",x"ca"),
   788 => (x"c4",x"49",x"f9",x"dc"),
   789 => (x"87",x"c4",x"86",x"70"),
   790 => (x"98",x"02",x"c1",x"f8"),
   791 => (x"87",x"c1",x"ca",x"c8"),
   792 => (x"bf",x"49",x"c7",x"ff"),
   793 => (x"81",x"c9",x"29",x"71"),
   794 => (x"7e",x"c0",x"4d",x"4c"),
   795 => (x"6e",x"48",x"c0",x"b7"),
   796 => (x"a8",x"06",x"c1",x"ef"),
   797 => (x"87",x"c1",x"c9",x"e0"),
   798 => (x"bf",x"49",x"c1",x"ca"),
   799 => (x"cc",x"bf",x"4a",x"c2"),
   800 => (x"8a",x"c1",x"c9",x"d0"),
   801 => (x"bf",x"4b",x"92",x"72"),
   802 => (x"a1",x"49",x"74",x"4a"),
   803 => (x"c1",x"c9",x"d4",x"bf"),
   804 => (x"9a",x"72",x"a1",x"49"),
   805 => (x"d4",x"66",x"1e",x"71"),
   806 => (x"e2",x"e6",x"87",x"c4"),
   807 => (x"86",x"70",x"98",x"05"),
   808 => (x"c5",x"87",x"c0",x"48"),
   809 => (x"c1",x"c2",x"87",x"c1"),
   810 => (x"84",x"74",x"49",x"c1"),
   811 => (x"c9",x"d4",x"bf",x"99"),
   812 => (x"05",x"ce",x"87",x"c1"),
   813 => (x"ca",x"cc",x"bf",x"49"),
   814 => (x"f5",x"f2",x"87",x"70"),
   815 => (x"49",x"c1",x"ca",x"d0"),
   816 => (x"59",x"d4",x"66",x"48"),
   817 => (x"c8",x"c0",x"80",x"d8"),
   818 => (x"a6",x"58",x"c1",x"85"),
   819 => (x"6e",x"b7",x"ad",x"04"),
   820 => (x"fe",x"e2",x"87",x"cf"),
   821 => (x"87",x"73",x"1e",x"c0"),
   822 => (x"f3",x"ed",x"1e",x"cb"),
   823 => (x"cf",x"87",x"c8",x"86"),
   824 => (x"c0",x"48",x"c5",x"87"),
   825 => (x"c1",x"ca",x"c8",x"bf"),
   826 => (x"48",x"26",x"e5",x"db"),
   827 => (x"87",x"43",x"61",x"6e"),
   828 => (x"27",x"74",x"20",x"6f"),
   829 => (x"70",x"65",x"6e",x"20"),
   830 => (x"25",x"73",x"0a",x"00"),
   831 => (x"1e",x"f3",x"48",x"71"),
   832 => (x"50",x"48",x"26",x"4f"),
   833 => (x"0e",x"5e",x"5b",x"5c"),
   834 => (x"5d",x"0e",x"f8",x"86"),
   835 => (x"71",x"4c",x"c0",x"e4"),
   836 => (x"66",x"4d",x"d5",x"fb"),
   837 => (x"a7",x"4b",x"c2",x"ca"),
   838 => (x"a7",x"7e",x"c4",x"a6"),
   839 => (x"48",x"c0",x"78",x"74"),
   840 => (x"9c",x"05",x"c6",x"87"),
   841 => (x"c0",x"f0",x"53",x"c1"),
   842 => (x"c6",x"87",x"74",x"9c"),
   843 => (x"02",x"c0",x"e2",x"87"),
   844 => (x"74",x"49",x"1e",x"dc"),
   845 => (x"66",x"4a",x"ca",x"ec"),
   846 => (x"87",x"71",x"4a",x"26"),
   847 => (x"49",x"6e",x"82",x"12"),
   848 => (x"53",x"d8",x"66",x"4a"),
   849 => (x"ca",x"de",x"87",x"70"),
   850 => (x"49",x"4c",x"c1",x"8d"),
   851 => (x"74",x"9c",x"05",x"ff"),
   852 => (x"de",x"87",x"c0",x"b7"),
   853 => (x"ad",x"06",x"d8",x"87"),
   854 => (x"c0",x"e8",x"66",x"02"),
   855 => (x"c5",x"87",x"c0",x"f0"),
   856 => (x"4a",x"c3",x"87",x"c0"),
   857 => (x"e0",x"4a",x"72",x"53"),
   858 => (x"c1",x"8d",x"c0",x"b7"),
   859 => (x"ad",x"01",x"e8",x"87"),
   860 => (x"d4",x"dd",x"a7",x"ab"),
   861 => (x"02",x"df",x"87",x"dc"),
   862 => (x"66",x"4c",x"c0",x"e0"),
   863 => (x"66",x"1e",x"c1",x"8b"),
   864 => (x"97",x"6b",x"49",x"74"),
   865 => (x"0f",x"c4",x"86",x"66"),
   866 => (x"48",x"c1",x"80",x"c8"),
   867 => (x"a6",x"58",x"d3",x"ff"),
   868 => (x"a7",x"ab",x"05",x"ff"),
   869 => (x"e4",x"87",x"c4",x"66"),
   870 => (x"48",x"f8",x"8e",x"26"),
   871 => (x"4d",x"26",x"4c",x"26"),
   872 => (x"4b",x"26",x"4f",x"30"),
   873 => (x"31",x"32",x"33",x"34"),
   874 => (x"35",x"36",x"37",x"38"),
   875 => (x"39",x"41",x"42",x"43"),
   876 => (x"44",x"45",x"46",x"00"),
   877 => (x"0e",x"5e",x"5b",x"5c"),
   878 => (x"5d",x"0e",x"71",x"4b"),
   879 => (x"ff",x"4d",x"13",x"4c"),
   880 => (x"9c",x"02",x"d7",x"87"),
   881 => (x"c1",x"85",x"d4",x"66"),
   882 => (x"1e",x"74",x"49",x"d4"),
   883 => (x"66",x"0f",x"c4",x"86"),
   884 => (x"74",x"a8",x"05",x"c6"),
   885 => (x"87",x"13",x"4c",x"9c"),
   886 => (x"05",x"e9",x"87",x"75"),
   887 => (x"48",x"26",x"4d",x"26"),
   888 => (x"4c",x"26",x"4b",x"26"),
   889 => (x"4f",x"0e",x"5e",x"5b"),
   890 => (x"5c",x"5d",x"0e",x"e8"),
   891 => (x"86",x"c8",x"a6",x"59"),
   892 => (x"c0",x"e8",x"66",x"4d"),
   893 => (x"c0",x"4c",x"c8",x"a6"),
   894 => (x"48",x"c0",x"78",x"c4"),
   895 => (x"66",x"97",x"bf",x"4b"),
   896 => (x"c4",x"66",x"48",x"c1"),
   897 => (x"80",x"c8",x"a6",x"58"),
   898 => (x"73",x"9b",x"02",x"c6"),
   899 => (x"d3",x"87",x"c8",x"66"),
   900 => (x"02",x"c5",x"d9",x"87"),
   901 => (x"cc",x"a6",x"48",x"c0"),
   902 => (x"78",x"fc",x"80",x"c0"),
   903 => (x"78",x"73",x"4a",x"c0"),
   904 => (x"e0",x"8a",x"02",x"c3"),
   905 => (x"c8",x"87",x"c3",x"8a"),
   906 => (x"02",x"c3",x"c2",x"87"),
   907 => (x"c2",x"8a",x"02",x"c2"),
   908 => (x"ea",x"87",x"8a",x"02"),
   909 => (x"c2",x"f7",x"87",x"c4"),
   910 => (x"8a",x"02",x"c2",x"f1"),
   911 => (x"87",x"c2",x"8a",x"02"),
   912 => (x"c2",x"eb",x"87",x"c3"),
   913 => (x"8a",x"02",x"c2",x"ed"),
   914 => (x"87",x"d4",x"8a",x"02"),
   915 => (x"c0",x"fa",x"87",x"8a"),
   916 => (x"02",x"c1",x"c5",x"87"),
   917 => (x"ca",x"8a",x"02",x"c0"),
   918 => (x"f7",x"87",x"c1",x"8a"),
   919 => (x"02",x"c1",x"e5",x"87"),
   920 => (x"8a",x"02",x"c0",x"e4"),
   921 => (x"87",x"c5",x"8a",x"02"),
   922 => (x"df",x"87",x"c3",x"8a"),
   923 => (x"02",x"c1",x"cd",x"87"),
   924 => (x"c4",x"8a",x"02",x"c0"),
   925 => (x"e3",x"87",x"c3",x"8a"),
   926 => (x"02",x"c0",x"e5",x"87"),
   927 => (x"c2",x"8a",x"02",x"c8"),
   928 => (x"87",x"c3",x"8a",x"02"),
   929 => (x"d3",x"87",x"c1",x"f9"),
   930 => (x"87",x"cc",x"a6",x"48"),
   931 => (x"ca",x"78",x"c2",x"d2"),
   932 => (x"87",x"cc",x"a6",x"48"),
   933 => (x"c2",x"78",x"c2",x"ca"),
   934 => (x"87",x"cc",x"a6",x"48"),
   935 => (x"d0",x"78",x"c2",x"c2"),
   936 => (x"87",x"c0",x"f0",x"66"),
   937 => (x"1e",x"c0",x"f0",x"66"),
   938 => (x"1e",x"c4",x"85",x"75"),
   939 => (x"4a",x"c4",x"8a",x"6a"),
   940 => (x"49",x"fc",x"c0",x"87"),
   941 => (x"c8",x"86",x"70",x"49"),
   942 => (x"a4",x"4c",x"c1",x"e6"),
   943 => (x"87",x"c8",x"a6",x"48"),
   944 => (x"c1",x"78",x"c1",x"de"),
   945 => (x"87",x"c0",x"f0",x"66"),
   946 => (x"1e",x"c4",x"85",x"75"),
   947 => (x"4a",x"c4",x"8a",x"6a"),
   948 => (x"49",x"c0",x"f0",x"66"),
   949 => (x"0f",x"c4",x"86",x"c1"),
   950 => (x"84",x"c1",x"c7",x"87"),
   951 => (x"c0",x"f0",x"66",x"1e"),
   952 => (x"c0",x"e5",x"49",x"c0"),
   953 => (x"f0",x"66",x"0f",x"c4"),
   954 => (x"86",x"c1",x"84",x"c0"),
   955 => (x"f5",x"87",x"c8",x"a6"),
   956 => (x"48",x"c1",x"78",x"c0"),
   957 => (x"ed",x"87",x"d0",x"a6"),
   958 => (x"48",x"c1",x"78",x"f8"),
   959 => (x"80",x"c1",x"78",x"c0"),
   960 => (x"e1",x"87",x"c0",x"f0"),
   961 => (x"ab",x"06",x"db",x"87"),
   962 => (x"c0",x"f9",x"ab",x"03"),
   963 => (x"d5",x"87",x"d4",x"66"),
   964 => (x"4a",x"ca",x"92",x"73"),
   965 => (x"49",x"c0",x"f0",x"89"),
   966 => (x"72",x"a1",x"49",x"d8"),
   967 => (x"a6",x"59",x"48",x"f4"),
   968 => (x"80",x"c1",x"78",x"cc"),
   969 => (x"66",x"02",x"c1",x"e5"),
   970 => (x"87",x"c4",x"85",x"75"),
   971 => (x"49",x"c4",x"89",x"69"),
   972 => (x"7e",x"c1",x"e4",x"ab"),
   973 => (x"05",x"d5",x"87",x"6e"),
   974 => (x"48",x"c0",x"b7",x"a8"),
   975 => (x"03",x"cd",x"87",x"c0"),
   976 => (x"ed",x"49",x"f6",x"f7"),
   977 => (x"87",x"6e",x"48",x"c0"),
   978 => (x"08",x"88",x"70",x"7e"),
   979 => (x"d0",x"66",x"1e",x"d8"),
   980 => (x"66",x"1e",x"c0",x"f8"),
   981 => (x"66",x"1e",x"c0",x"f8"),
   982 => (x"66",x"1e",x"dc",x"66"),
   983 => (x"49",x"1e",x"d4",x"66"),
   984 => (x"49",x"f6",x"e0",x"87"),
   985 => (x"d4",x"86",x"70",x"49"),
   986 => (x"a4",x"4c",x"c0",x"e1"),
   987 => (x"87",x"c0",x"e5",x"ab"),
   988 => (x"05",x"cf",x"87",x"d0"),
   989 => (x"a6",x"48",x"c0",x"78"),
   990 => (x"c4",x"80",x"c0",x"78"),
   991 => (x"f4",x"80",x"c1",x"78"),
   992 => (x"cc",x"87",x"c0",x"f0"),
   993 => (x"66",x"1e",x"73",x"49"),
   994 => (x"c0",x"f0",x"66",x"0f"),
   995 => (x"c4",x"86",x"c4",x"66"),
   996 => (x"97",x"bf",x"4b",x"c4"),
   997 => (x"66",x"48",x"c1",x"80"),
   998 => (x"c8",x"a6",x"58",x"73"),
   999 => (x"9b",x"05",x"f9",x"ed"),
  1000 => (x"87",x"74",x"48",x"e8"),
  1001 => (x"8e",x"26",x"4d",x"26"),
  1002 => (x"4c",x"26",x"4b",x"26"),
  1003 => (x"4f",x"1e",x"c0",x"1e"),
  1004 => (x"f5",x"c9",x"a7",x"1e"),
  1005 => (x"d0",x"a6",x"1e",x"d0"),
  1006 => (x"66",x"49",x"f8",x"e8"),
  1007 => (x"87",x"f4",x"8e",x"26"),
  1008 => (x"4f",x"0e",x"5e",x"5b"),
  1009 => (x"5c",x"0e",x"71",x"4b"),
  1010 => (x"c0",x"4c",x"13",x"4a"),
  1011 => (x"9a",x"02",x"cd",x"87"),
  1012 => (x"72",x"49",x"f4",x"e7"),
  1013 => (x"87",x"c1",x"84",x"13"),
  1014 => (x"4a",x"9a",x"05",x"f3"),
  1015 => (x"87",x"74",x"48",x"26"),
  1016 => (x"4c",x"26",x"4b",x"26"),
  1017 => (x"4f",x"1e",x"73",x"1e"),
  1018 => (x"72",x"9a",x"02",x"c0"),
  1019 => (x"e7",x"87",x"c0",x"48"),
  1020 => (x"c1",x"4b",x"72",x"a9"),
  1021 => (x"06",x"d1",x"87",x"72"),
  1022 => (x"82",x"06",x"c9",x"87"),
  1023 => (x"73",x"83",x"72",x"a9"),
  1024 => (x"01",x"f4",x"87",x"c3"),
  1025 => (x"87",x"c1",x"b2",x"3a"),
  1026 => (x"72",x"a9",x"03",x"89"),
  1027 => (x"73",x"80",x"07",x"c1"),
  1028 => (x"2a",x"2b",x"05",x"f3"),
  1029 => (x"87",x"26",x"4b",x"26"),
  1030 => (x"4f",x"1e",x"75",x"1e"),
  1031 => (x"c4",x"4d",x"71",x"b7"),
  1032 => (x"a1",x"04",x"ff",x"b9"),
  1033 => (x"c1",x"81",x"c3",x"bd"),
  1034 => (x"07",x"72",x"b7",x"a2"),
  1035 => (x"04",x"ff",x"ba",x"c1"),
  1036 => (x"82",x"c1",x"bd",x"07"),
  1037 => (x"fe",x"ee",x"87",x"c1"),
  1038 => (x"2d",x"04",x"ff",x"b8"),
  1039 => (x"c1",x"80",x"07",x"2d"),
  1040 => (x"04",x"ff",x"b9",x"c1"),
  1041 => (x"81",x"07",x"26",x"4d"),
  1042 => (x"26",x"4f",x"26",x"4d"),
	others => (others => x"00")
);

-- Xilinx XST attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "no_rw_check";

-- Altera Quartus attributes
attribute ramstyle: string;
attribute ramstyle of ram: signal is "no_rw_check";

signal q_local : word_t;
signal q2_local : word_t;

begin
    
	process(clk,q_local)
	begin

		q(31 downto 24)<=q_local(0);
		q(23 downto 16)<=q_local(1);
		q(15 downto 8)<=q_local(2);
		q(7 downto 0)<=q_local(3);

		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel(3) = '1') then
					ram(to_integer(unsigned(addr)))(3) <= d(7 downto 0);
				end if;
				if bytesel(2) = '1' then
					ram(to_integer(unsigned(addr)))(2) <= d(15 downto 8);
				end if;
				if bytesel(1) = '1' then
					ram(to_integer(unsigned(addr)))(1) <= d(23 downto 16);
				end if;
				if bytesel(0) = '1' then
					ram(to_integer(unsigned(addr)))(0) <= d(31 downto 24);
				end if;
			end if;
			q_local <= ram(to_integer(unsigned(addr)));
		end if;
	end process;

	-- Second port
	
	process(clk,q2_local)
	begin

		q2(31 downto 24)<=q2_local(0);
		q2(23 downto 16)<=q2_local(1);
		q2(15 downto 8)<=q2_local(2);
		q2(7 downto 0)<=q2_local(3);

		if(rising_edge(clk)) then 
			if(we2 = '1') then
				-- edit this code if using other than four bytes per word
				if(bytesel2(3) = '1') then
					ram(to_integer(unsigned(addr2)))(3) <= d2(7 downto 0);
				end if;
				if bytesel2(2) = '1' then
					ram(to_integer(unsigned(addr2)))(2) <= d2(15 downto 8);
				end if;
				if bytesel2(1) = '1' then
					ram(to_integer(unsigned(addr2)))(1) <= d2(23 downto 16);
				end if;
				if bytesel2(0) = '1' then
					ram(to_integer(unsigned(addr2)))(0) <= d2(31 downto 24);
				end if;
			end if;
			q2_local <= ram(to_integer(unsigned(addr2)));
		end if;
	end process;

end arch;

